#supernode.ckt
.circuit
Vsource1 2 3  dc 22
I1 1 2 dc 3
I2 1 GND DC 8
I3 GND 3 DC 25
R1 1 3 4
R2 1 2 3
R3 2 GND 1 
R4 3 GND 5
.end
